dmel OreR F AC R1 201883 81407 138509
dmel OreR F AC R2 193274 72883 105452
dmel OreR F AC R3 216127 85068 136064
dmel OreR F AC R4 261609 114350 179157
dmel OreR F GO R1 24858 8839 37701
dmel OreR F GO R2 19485 8434 34577
dmel OreR F GO R3 9519 4652 16701
dmel OreR F GO R4 13553 6259 21778
dmel OreR F HD R1 200120 96002 143413
dmel OreR F HD R2 170495 82897 106357
dmel OreR F HD R3 205158 116974 130450
dmel OreR F HD R4 235198 113107 165446
dmel OreR F IR R1 242928 104052 151759
dmel OreR F IR R2 223021 97050 127410
dmel OreR F IR R3 195422 80660 117279
dmel OreR F IR R4 257440 126931 168682
dmel OreR F TE R1 17055 6539 10035
dmel OreR F TE R2 76164 26756 38099
dmel OreR F TE R3 20465 8869 12840
dmel OreR F TE R4 72228 32505 47613
dmel OreR F TX R1 124298 60049 88435
dmel OreR F TX R2 110510 52932 66480
dmel OreR F TX R3 125785 70679 79639
dmel OreR F TX R4 150159 85050 102885
dmel OreR F VS R1 10851 4910 7695
dmel OreR F VS R2 4187 1908 2563
dmel OreR F VS R3 6440 2559 4057
dmel OreR F VS R4 5290 2494 3792
dmel OreR F WO R1 102602 37509 81493
dmel OreR F WO R2 61021 28563 54461
dmel OreR F WO R3 58254 25225 43341
dmel OreR F WO R4 96194 47126 82891
dmel OreR M AC R1 34 28 27
dmel OreR M AC R2 44 20 21
dmel OreR M AC R3 69 45 62
dmel OreR M AC R4 61 69 57
dmel OreR M GO R1 11 7 8
dmel OreR M GO R2 90 60 73
dmel OreR M GO R3 30 19 38
dmel OreR M GO R4 29 18 27
dmel OreR M HD R1 71 68 53
dmel OreR M HD R2 42 137 37
dmel OreR M HD R3 61 106 64
dmel OreR M HD R4 76 117 65
dmel OreR M IR R1 42 26 30
dmel OreR M IR R2 1 2 1
dmel OreR M IR R3 42 28 36
dmel OreR M IR R4 147 42 76
dmel OreR M TE R1 52 36 24
dmel OreR M TE R2 7 3 5
dmel OreR M TE R3 2 4 2
dmel OreR M TE R4 210 93 128
dmel OreR M TX R1 18 33 11
dmel OreR M TX R2 33 24 38
dmel OreR M TX R3 52 49 43
dmel OreR M TX R4 32 36 32
dmel OreR M VS R1 3 11 1
dmel OreR M VS R2 3 14 3
dmel OreR M VS R3 4 12 2
dmel OreR M VS R4 2 19 2
dmel OreR M WO R1 12 18 11
dmel OreR M WO R2 44 30 58
dmel OreR M WO R3 2 38 5
dmel OreR M WO R4 30 37 44
dmel w1118 F AC R1 298361 137189 186157
dmel w1118 F AC R2 227868 92073 133473
dmel w1118 F AC R3 269822 116657 135688
dmel w1118 F AC R4 130360 59343 59072
dmel w1118 F GO R1 14126 10516 26050
dmel w1118 F GO R2 9570 7448 17521
dmel w1118 F GO R3 10271 9209 19640
dmel w1118 F GO R4 8057 7007 16415
dmel w1118 F HD R1 131881 105862 66269
dmel w1118 F HD R2 141101 83492 45443
dmel w1118 F HD R3 209026 154590 87596
dmel w1118 F HD R4 163010 114186 59865
dmel w1118 F IR R1 133552 59382 83971
dmel w1118 F IR R2 144879 69513 86276
dmel w1118 F IR R3 238121 116018 130595
dmel w1118 F IR R4 134394 70499 68996
dmel w1118 F TE R1 43220 19573 27063
dmel w1118 F TE R2 9418 4449 4956
dmel w1118 F TE R3 6969 3501 3215
dmel w1118 F TE R4 33735 14493 14322
dmel w1118 F TX R1 65490 51818 28623
dmel w1118 F TX R2 94643 62125 34664
dmel w1118 F TX R3 83276 63307 36359
dmel w1118 F TX R4 94721 79447 42135
dmel w1118 F VS R1 4740 2184 3285
dmel w1118 F VS R2 2734 1512 1772
dmel w1118 F VS R3 2292 1311 1420
dmel w1118 F VS R4 2094 1197 1044
dmel w1118 F WO R1 26511 15288 21316
dmel w1118 F WO R2 50394 26440 32956
dmel w1118 F WO R3 51220 28082 36008
dmel w1118 F WO R4 93948 36591 44902
dmel w1118 M AC R1 33 21 15
dmel w1118 M AC R2 1 1 5
dmel w1118 M AC R3 29 11 18
dmel w1118 M AC R4 34 26 32
dmel w1118 M GO R1 0 4 2
dmel w1118 M GO R2 3 2 3
dmel w1118 M GO R3 0 7 2
dmel w1118 M GO R4 0 7 7
dmel w1118 M HD R1 4 274 4
dmel w1118 M HD R2 49 356 22
dmel w1118 M HD R3 31 176 16
dmel w1118 M HD R4 89 331 25
dmel w1118 M IR R1 33 10 37
dmel w1118 M IR R2 32 19 17
dmel w1118 M IR R3 34 13 13
dmel w1118 M IR R4 5 3 2
dmel w1118 M TE R1 20 12 15
dmel w1118 M TE R2 2 3 1
dmel w1118 M TE R3 7 5 6
dmel w1118 M TE R4 2 0 2
dmel w1118 M TX R1 12 9 11
dmel w1118 M TX R2 9 12 8
dmel w1118 M TX R3 13 18 3
dmel w1118 M TX R4 28 22 8
dmel w1118 M VS R1 8 41 2
dmel w1118 M VS R2 1 36 1
dmel w1118 M VS R3 0 41 1
dmel w1118 M VS R4 0 53 3
dmel w1118 M WO R1 5 41 4
dmel w1118 M WO R2 1 38 10
dmel w1118 M WO R3 4 48 11
dmel w1118 M WO R4 5 38 6
